// timer_display_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module timer_display_tb (
	);

	wire         timer_display_inst_clk_bfm_clk_clk;                 // timer_display_inst_clk_bfm:clk -> [timer_display_inst:clk_clk, timer_display_inst_reset_bfm:clk]
	wire  [27:0] timer_display_inst_display_7_segments_export;       // timer_display_inst:display_7_segments_export -> timer_display_inst_display_7_segments_bfm:sig_export
	wire   [0:0] timer_display_inst_pause_button_bfm_conduit_export; // timer_display_inst_pause_button_bfm:sig_export -> timer_display_inst:pause_button_export
	wire   [0:0] timer_display_inst_reset_button_bfm_conduit_export; // timer_display_inst_reset_button_bfm:sig_export -> timer_display_inst:reset_button_export
	wire   [0:0] timer_display_inst_start_button_bfm_conduit_export; // timer_display_inst_start_button_bfm:sig_export -> timer_display_inst:start_button_export
	wire         timer_display_inst_reset_bfm_reset_reset;           // timer_display_inst_reset_bfm:reset -> timer_display_inst:reset_reset_n

	timer_display timer_display_inst (
		.clk_clk                   (timer_display_inst_clk_bfm_clk_clk),                 //                clk.clk
		.display_7_segments_export (timer_display_inst_display_7_segments_export),       // display_7_segments.export
		.pause_button_export       (timer_display_inst_pause_button_bfm_conduit_export), //       pause_button.export
		.reset_reset_n             (timer_display_inst_reset_bfm_reset_reset),           //              reset.reset_n
		.reset_button_export       (timer_display_inst_reset_button_bfm_conduit_export), //       reset_button.export
		.start_button_export       (timer_display_inst_start_button_bfm_conduit_export)  //       start_button.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) timer_display_inst_clk_bfm (
		.clk (timer_display_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm timer_display_inst_display_7_segments_bfm (
		.sig_export (timer_display_inst_display_7_segments_export)  // conduit.export
	);

	altera_conduit_bfm_0002 timer_display_inst_pause_button_bfm (
		.sig_export (timer_display_inst_pause_button_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) timer_display_inst_reset_bfm (
		.reset (timer_display_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (timer_display_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 timer_display_inst_reset_button_bfm (
		.sig_export (timer_display_inst_reset_button_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 timer_display_inst_start_button_bfm (
		.sig_export (timer_display_inst_start_button_bfm_conduit_export)  // conduit.export
	);

endmodule
